library verilog;
use verilog.vl_types.all;
entity song_reader_tb is
end song_reader_tb;
