library verilog;
use verilog.vl_types.all;
entity note_player_tb is
end note_player_tb;
