library verilog;
use verilog.vl_types.all;
entity wave_display_top_tb is
end wave_display_top_tb;
