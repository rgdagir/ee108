library verilog;
use verilog.vl_types.all;
entity mcu_tb is
end mcu_tb;
