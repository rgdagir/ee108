library verilog;
use verilog.vl_types.all;
entity music_player_tb is
end music_player_tb;
