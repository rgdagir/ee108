library verilog;
use verilog.vl_types.all;
entity sine_reader_tb is
end sine_reader_tb;
