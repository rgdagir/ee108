library verilog;
use verilog.vl_types.all;
entity wave_display_tb is
end wave_display_tb;
