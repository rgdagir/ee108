library verilog;
use verilog.vl_types.all;
entity wave_capture_tb is
end wave_capture_tb;
