/*
 * A simple fake RAM that you can use to aid in debugging your wave display.
 */
module fake_sample_ram (
    input clk,
    input [7:0] addr,
    output reg [7:0] dout
);
	 wire [19:0] memory [511:0];
    always @(posedge clk)
        dout = memory[addr];

 assign memory [9'd  0] = 8'b10101001; 
 assign memory [9'd  1] = 8'b11001100; 
 assign memory [9'd  2] = 8'b11100111; 
 assign memory [9'd  3] = 8'b11111001; 
 assign memory [9'd  4] = 8'b11111111; 
 assign memory [9'd  5] = 8'b11111010; 
 assign memory [9'd  6] = 8'b11101000; 
 assign memory [9'd  7] = 8'b11001101; 
 assign memory [9'd  8] = 8'b10101011; 
 assign memory [9'd  9] = 8'b10000100; 
 assign memory [9'd 10] = 8'b01011110; 
 assign memory [9'd 11] = 8'b00111010; 
 assign memory [9'd 12] = 8'b00011101; 
 assign memory [9'd 13] = 8'b00001001; 
 assign memory [9'd 14] = 8'b00000000; 
 assign memory [9'd 15] = 8'b00000011; 
 assign memory [9'd 16] = 8'b00010010; 
 assign memory [9'd 17] = 8'b00101011; 
 assign memory [9'd 18] = 8'b01001101; 
 assign memory [9'd 19] = 8'b01110011; 
 assign memory [9'd 20] = 8'b10011010; 
 assign memory [9'd 21] = 8'b10111110; 
 assign memory [9'd 22] = 8'b11011101; 
 assign memory [9'd 23] = 8'b11110011; 
 assign memory [9'd 24] = 8'b11111110; 
 assign memory [9'd 25] = 8'b11111110; 
 assign memory [9'd 26] = 8'b11110001; 
 assign memory [9'd 27] = 8'b11011001; 
 assign memory [9'd 28] = 8'b10111010; 
 assign memory [9'd 29] = 8'b10010100; 
 assign memory [9'd 30] = 8'b01101101; 
 assign memory [9'd 31] = 8'b01001000; 
 assign memory [9'd 32] = 8'b00101000; 
 assign memory [9'd 33] = 8'b00001111; 
 assign memory [9'd 34] = 8'b00000010; 
 assign memory [9'd 35] = 8'b00000000; 
 assign memory [9'd 36] = 8'b00001011; 
 assign memory [9'd 37] = 8'b00100000; 
 assign memory [9'd 38] = 8'b00111110; 
 assign memory [9'd 39] = 8'b01100011; 
 assign memory [9'd 40] = 8'b10001010; 
 assign memory [9'd 41] = 8'b10110000; 
 assign memory [9'd 42] = 8'b11010010; 
 assign memory [9'd 43] = 8'b11101011; 
 assign memory [9'd 44] = 8'b11111011; 
 assign memory [9'd 45] = 8'b11111111; 
 assign memory [9'd 46] = 8'b11110111; 
 assign memory [9'd 47] = 8'b11110110; 
 assign memory [9'd 48] = 8'b11110110; 
 assign memory [9'd 49] = 8'b11110101; 
 assign memory [9'd 50] = 8'b11110100; 
 assign memory [9'd 51] = 8'b11110011; 
 assign memory [9'd 52] = 8'b11110001; 
 assign memory [9'd 53] = 8'b11110000; 
 assign memory [9'd 54] = 8'b11101111; 
 assign memory [9'd 55] = 8'b11101110; 
 assign memory [9'd 56] = 8'b11101101; 
 assign memory [9'd 57] = 8'b11101011; 
 assign memory [9'd 58] = 8'b11101010; 
 assign memory [9'd 59] = 8'b11101001; 
 assign memory [9'd 60] = 8'b11100111; 
 assign memory [9'd 61] = 8'b11100110; 
 assign memory [9'd 62] = 8'b11100100; 
 assign memory [9'd 63] = 8'b11100011; 
 assign memory [9'd 64] = 8'b11100001; 
 assign memory [9'd 65] = 8'b11011111; 
 assign memory [9'd 66] = 8'b11011110; 
 assign memory [9'd 67] = 8'b11011100; 
 assign memory [9'd 68] = 8'b11011010; 
 assign memory [9'd 69] = 8'b11011001; 
 assign memory [9'd 70] = 8'b11010111; 
 assign memory [9'd 71] = 8'b11010101; 
 assign memory [9'd 72] = 8'b11010011; 
 assign memory [9'd 73] = 8'b11010001; 
 assign memory [9'd 74] = 8'b11001111; 
 assign memory [9'd 75] = 8'b11001101; 
 assign memory [9'd 76] = 8'b11001011; 
 assign memory [9'd 77] = 8'b11001010; 
 assign memory [9'd 78] = 8'b11000111; 
 assign memory [9'd 79] = 8'b11000101; 
 assign memory [9'd 80] = 8'b11000011; 
 assign memory [9'd 81] = 8'b11000001; 
 assign memory [9'd 82] = 8'b10011000; 
 assign memory [9'd 83] = 8'b01101100; 
 assign memory [9'd 84] = 8'b01000011; 
 assign memory [9'd 85] = 8'b00100000; 
 assign memory [9'd 86] = 8'b00001001; 
 assign memory [9'd 88] = 8'b00000110; 
 assign memory [9'd 89] = 8'b00011010; 
 assign memory [9'd 90] = 8'b00111010; 
 assign memory [9'd 91] = 8'b01100011; 
 assign memory [9'd 92] = 8'b10001111; 
 assign memory [9'd 93] = 8'b10111001; 
 assign memory [9'd 94] = 8'b11011100; 
 assign memory [9'd 95] = 8'b11110101; 
 assign memory [9'd 96] = 8'b11111111; 
 assign memory [9'd 97] = 8'b11111011; 
 assign memory [9'd 98] = 8'b11100111; 
 assign memory [9'd 99] = 8'b11001000; 
 assign memory [9'd100] = 8'b10100000; 
 assign memory [9'd101] = 8'b01110100; 
 assign memory [9'd102] = 8'b01001010; 
 assign memory [9'd103] = 8'b00100110; 
 assign memory [9'd104] = 8'b00001100; 
 assign memory [9'd105] = 8'b00000000; 
 assign memory [9'd106] = 8'b00000011; 
 assign memory [9'd107] = 8'b00010101; 
 assign memory [9'd108] = 8'b00110100; 
 assign memory [9'd109] = 8'b01011011; 
 assign memory [9'd110] = 8'b10000111; 
 assign memory [9'd111] = 8'b10110010; 
 assign memory [9'd112] = 8'b11010110; 
 assign memory [9'd113] = 8'b11110001; 
 assign memory [9'd114] = 8'b11111110; 
 assign memory [9'd115] = 8'b11111101; 
 assign memory [9'd116] = 8'b11101100; 
 assign memory [9'd117] = 8'b11001111; 
 assign memory [9'd118] = 8'b10101000; 
 assign memory [9'd119] = 8'b01111100; 
 assign memory [9'd120] = 8'b01010001; 
 assign memory [9'd121] = 8'b00101011; 
 assign memory [9'd122] = 8'b00010000; 
 assign memory [9'd123] = 8'b00000001; 
 assign memory [9'd124] = 8'b00000010; 
 assign memory [9'd125] = 8'b00010001; 
 assign memory [9'd126] = 8'b00101101; 
 assign memory [9'd127] = 8'b01010011; 
 assign memory [9'd128] = 8'b01111111; 
 assign memory [9'd129] = 8'b10101010; 
 assign memory [9'd130] = 8'b11010000; 
 assign memory [9'd131] = 8'b11101101; 
 assign memory [9'd132] = 8'b11111101; 
 assign memory [9'd133] = 8'b11111110; 
 assign memory [9'd134] = 8'b11110000; 
 assign memory [9'd135] = 8'b11101111; 
 assign memory [9'd136] = 8'b11101101; 
 assign memory [9'd137] = 8'b11101100; 
 assign memory [9'd139] = 8'b11101001; 
 assign memory [9'd140] = 8'b11100111; 
 assign memory [9'd141] = 8'b11100101; 
 assign memory [9'd142] = 8'b11100100; 
 assign memory [9'd143] = 8'b11100010; 
 assign memory [9'd144] = 8'b11100000; 
 assign memory [9'd145] = 8'b11011110; 
 assign memory [9'd146] = 8'b11011101; 
 assign memory [9'd147] = 8'b11011011; 
 assign memory [9'd148] = 8'b11011001; 
 assign memory [9'd149] = 8'b11010111; 
 assign memory [9'd150] = 8'b11010101; 
 assign memory [9'd151] = 8'b11010011; 
 assign memory [9'd152] = 8'b11010000; 
 assign memory [9'd153] = 8'b11001110; 
 assign memory [9'd154] = 8'b11001100; 
 assign memory [9'd155] = 8'b11001010; 
 assign memory [9'd156] = 8'b11001000; 
 assign memory [9'd157] = 8'b11000101; 
 assign memory [9'd158] = 8'b11000011; 
 assign memory [9'd159] = 8'b11000001; 
 assign memory [9'd160] = 8'b10111110; 
 assign memory [9'd161] = 8'b10111100; 
 assign memory [9'd162] = 8'b10111001; 
 assign memory [9'd163] = 8'b10110111; 
 assign memory [9'd164] = 8'b10110100; 
 assign memory [9'd165] = 8'b10110010; 
 assign memory [9'd166] = 8'b10101111; 
 assign memory [9'd167] = 8'b10101101; 
 assign memory [9'd168] = 8'b10101010; 
 assign memory [9'd169] = 8'b10100111; 
 assign memory [9'd170] = 8'b01111010; 
 assign memory [9'd171] = 8'b01001100; 
 assign memory [9'd172] = 8'b00100110; 
 assign memory [9'd173] = 8'b00001011; 
 assign memory [9'd174] = 8'b00000000; 
 assign memory [9'd175] = 8'b00000101; 
 assign memory [9'd176] = 8'b00011011; 
 assign memory [9'd177] = 8'b00111110; 
 assign memory [9'd178] = 8'b01101010; 
 assign memory [9'd179] = 8'b10011000; 
 assign memory [9'd180] = 8'b11000011; 
 assign memory [9'd181] = 8'b11100110; 
 assign memory [9'd182] = 8'b11111010; 
 assign memory [9'd183] = 8'b11111111; 
 assign memory [9'd184] = 8'b11110011; 
 assign memory [9'd185] = 8'b11010111; 
 assign memory [9'd186] = 8'b10110000; 
 assign memory [9'd187] = 8'b10000010; 
 assign memory [9'd188] = 8'b01010101; 
 assign memory [9'd189] = 8'b00101100; 
 assign memory [9'd190] = 8'b00001111; 
 assign memory [9'd191] = 8'b00000001; 
 assign memory [9'd192] = 8'b00000011; 
 assign memory [9'd193] = 8'b00010110; 
 assign memory [9'd194] = 8'b00110111; 
 assign memory [9'd195] = 8'b01100001; 
 assign memory [9'd196] = 8'b10001111; 
 assign memory [9'd197] = 8'b10111100; 
 assign memory [9'd198] = 8'b11100000; 
 assign memory [9'd199] = 8'b11111000; 
 assign memory [9'd200] = 8'b11111111; 
 assign memory [9'd201] = 8'b11110110; 
 assign memory [9'd202] = 8'b11011101; 
 assign memory [9'd203] = 8'b10111000; 
 assign memory [9'd204] = 8'b10001011; 
 assign memory [9'd205] = 8'b01011101; 
 assign memory [9'd206] = 8'b00110011; 
 assign memory [9'd207] = 8'b00010100; 
 assign memory [9'd208] = 8'b00000010; 
 assign memory [9'd209] = 8'b00000001; 
 assign memory [9'd210] = 8'b00010001; 
 assign memory [9'd211] = 8'b00101111; 
 assign memory [9'd212] = 8'b01011000; 
 assign memory [9'd213] = 8'b10000110; 
 assign memory [9'd214] = 8'b10110100; 
 assign memory [9'd215] = 8'b11011010; 
 assign memory [9'd216] = 8'b11110100; 
 assign memory [9'd217] = 8'b11111111; 
 assign memory [9'd218] = 8'b11111001; 
 assign memory [9'd219] = 8'b11100011; 
 assign memory [9'd220] = 8'b11000000; 
 assign memory [9'd221] = 8'b10010100; 
 assign memory [9'd222] = 8'b01100110; 
 assign memory [9'd223] = 8'b01100011; 
 assign memory [9'd224] = 8'b01100000; 
 assign memory [9'd225] = 8'b01011101; 
 assign memory [9'd226] = 8'b01011011; 
 assign memory [9'd227] = 8'b01011000; 
 assign memory [9'd228] = 8'b01010101; 
 assign memory [9'd229] = 8'b01010010; 
 assign memory [9'd230] = 8'b01010000; 
 assign memory [9'd231] = 8'b01001101; 
 assign memory [9'd232] = 8'b01001010; 
 assign memory [9'd233] = 8'b01001000; 
 assign memory [9'd234] = 8'b01000101; 
 assign memory [9'd235] = 8'b01000010; 
 assign memory [9'd236] = 8'b01000000; 
 assign memory [9'd237] = 8'b00111101; 
 assign memory [9'd238] = 8'b00111011; 
 assign memory [9'd239] = 8'b00111000; 
 assign memory [9'd240] = 8'b00110110; 
 assign memory [9'd241] = 8'b00110100; 
 assign memory [9'd242] = 8'b00110001; 
 assign memory [9'd243] = 8'b00101111; 
 assign memory [9'd244] = 8'b00101101; 
 assign memory [9'd245] = 8'b00101010; 
 assign memory [9'd246] = 8'b00101000; 
 assign memory [9'd247] = 8'b00100110; 
 assign memory [9'd248] = 8'b00100100; 
 assign memory [9'd249] = 8'b00100010; 
 assign memory [9'd250] = 8'b00100000; 
 assign memory [9'd251] = 8'b00011110; 
 assign memory [9'd252] = 8'b00011100; 
 assign memory [9'd253] = 8'b00011010; 
 assign memory [9'd254] = 8'b00011001; 
 assign memory [9'd255] = 8'b00010111; 
 assign memory [9'd256] = 8'b11010101; 
 assign memory [9'd257] = 8'b11110100; 
 assign memory [9'd258] = 8'b11111111; 
 assign memory [9'd259] = 8'b11110110; 
 assign memory [9'd260] = 8'b11011000; 
 assign memory [9'd261] = 8'b10101100; 
 assign memory [9'd262] = 8'b01111001; 
 assign memory [9'd263] = 8'b01000110; 
 assign memory [9'd264] = 8'b00011101; 
 assign memory [9'd265] = 8'b00000101; 
 assign memory [9'd266] = 8'b00000001; 
 assign memory [9'd267] = 8'b00010010; 
 assign memory [9'd268] = 8'b00110101; 
 assign memory [9'd269] = 8'b01100100; 
 assign memory [9'd270] = 8'b10011000; 
 assign memory [9'd271] = 8'b11001001; 
 assign memory [9'd272] = 8'b11101100; 
 assign memory [9'd273] = 8'b11111110; 
 assign memory [9'd274] = 8'b11111011; 
 assign memory [9'd275] = 8'b11100011; 
 assign memory [9'd276] = 8'b10111011; 
 assign memory [9'd277] = 8'b10001001; 
 assign memory [9'd278] = 8'b01010101; 
 assign memory [9'd279] = 8'b00101000; 
 assign memory [9'd280] = 8'b00001010; 
 assign memory [9'd281] = 8'b00000000; 
 assign memory [9'd282] = 8'b00001010; 
 assign memory [9'd283] = 8'b00101000; 
 assign memory [9'd284] = 8'b01010101; 
 assign memory [9'd285] = 8'b10001001; 
 assign memory [9'd286] = 8'b10111011; 
 assign memory [9'd287] = 8'b11100011; 
 assign memory [9'd288] = 8'b11111011; 
 assign memory [9'd289] = 8'b11111110; 
 assign memory [9'd290] = 8'b11101100; 
 assign memory [9'd291] = 8'b11001000; 
 assign memory [9'd292] = 8'b10011000; 
 assign memory [9'd293] = 8'b01100100; 
 assign memory [9'd294] = 8'b00110101; 
 assign memory [9'd295] = 8'b00010010; 
 assign memory [9'd296] = 8'b00000001; 
 assign memory [9'd297] = 8'b00000101; 
 assign memory [9'd298] = 8'b00011101; 
 assign memory [9'd299] = 8'b01000110; 
 assign memory [9'd300] = 8'b01111001; 
 assign memory [9'd301] = 8'b10101100; 
 assign memory [9'd302] = 8'b11011000; 
 assign memory [9'd303] = 8'b11011011; 
 assign memory [9'd304] = 8'b11011101; 
 assign memory [9'd305] = 8'b11011111; 
 assign memory [9'd306] = 8'b11100001; 
 assign memory [9'd307] = 8'b11100011; 
 assign memory [9'd308] = 8'b11100101; 
 assign memory [9'd309] = 8'b11100111; 
 assign memory [9'd310] = 8'b11101001; 
 assign memory [9'd311] = 8'b11101011; 
 assign memory [9'd312] = 8'b11101101; 
 assign memory [9'd313] = 8'b11101110; 
 assign memory [9'd314] = 8'b11110000; 
 assign memory [9'd315] = 8'b11110010; 
 assign memory [9'd316] = 8'b11110011; 
 assign memory [9'd317] = 8'b11110100; 
 assign memory [9'd318] = 8'b11110110; 
 assign memory [9'd319] = 8'b11110111; 
 assign memory [9'd320] = 8'b11111000; 
 assign memory [9'd321] = 8'b11111001; 
 assign memory [9'd322] = 8'b11111010; 
 assign memory [9'd323] = 8'b11111011; 
 assign memory [9'd324] = 8'b11111100; 
 assign memory [9'd325] = 8'b11111101; 
 assign memory [9'd326] = 8'b11111101; 
 assign memory [9'd327] = 8'b11111110; 
 assign memory [9'd328] = 8'b11111110; 
 assign memory [9'd329] = 8'b11111111; 
 assign memory [9'd330] = 8'b11111111; 
 assign memory [9'd331] = 8'b11111111; 
 assign memory [9'd332] = 8'b11111111; 
 assign memory [9'd333] = 8'b11111111; 
 assign memory [9'd334] = 8'b11111111; 
 assign memory [9'd335] = 8'b11111111; 
 assign memory [9'd336] = 8'b11111111; 
 assign memory [9'd337] = 8'b11111111; 
 assign memory [9'd338] = 8'b11111111; 
 assign memory [9'd339] = 8'b11111110; 
 assign memory [9'd340] = 8'b11111101; 
 assign memory [9'd341] = 8'b11111101; 
 assign memory [9'd342] = 8'b11111100; 
 assign memory [9'd343] = 8'b11111011; 
 assign memory [9'd344] = 8'b11111010; 
 assign memory [9'd345] = 8'b11111001; 
 assign memory [9'd346] = 8'b11111000; 
 assign memory [9'd347] = 8'b11110110; 
 assign memory [9'd348] = 8'b11110101; 
 assign memory [9'd349] = 8'b11110011; 
 assign memory [9'd350] = 8'b11110010; 
 assign memory [9'd351] = 8'b11110000; 
 assign memory [9'd352] = 8'b11101110; 
 assign memory [9'd353] = 8'b11101100; 
 assign memory [9'd354] = 8'b11101010; 
 assign memory [9'd355] = 8'b11101000; 
 assign memory [9'd356] = 8'b11100110; 
 assign memory [9'd357] = 8'b11100100; 
 assign memory [9'd358] = 8'b11100001; 
 assign memory [9'd359] = 8'b11011111; 
 assign memory [9'd360] = 8'b11011100; 
 assign memory [9'd361] = 8'b11011010; 
 assign memory [9'd362] = 8'b11010111; 
 assign memory [9'd363] = 8'b11010101; 
 assign memory [9'd364] = 8'b11010010; 
 assign memory [9'd365] = 8'b11001111; 
 assign memory [9'd366] = 8'b11001100; 
 assign memory [9'd367] = 8'b11001001; 
 assign memory [9'd368] = 8'b11000110; 
 assign memory [9'd369] = 8'b11000011; 
 assign memory [9'd370] = 8'b11000000; 
 assign memory [9'd371] = 8'b10111101; 
 assign memory [9'd372] = 8'b10111001; 
 assign memory [9'd373] = 8'b10110110; 
 assign memory [9'd374] = 8'b10110011; 
 assign memory [9'd375] = 8'b10101111; 
 assign memory [9'd376] = 8'b10101100; 
 assign memory [9'd377] = 8'b10101000; 
 assign memory [9'd378] = 8'b10100101; 
 assign memory [9'd379] = 8'b10100001; 
 assign memory [9'd380] = 8'b10011110; 
 assign memory [9'd381] = 8'b10011010; 
 assign memory [9'd382] = 8'b10010110; 
 assign memory [9'd383] = 8'b10010011; 
 assign memory [9'd384] = 8'b10001111; 
 assign memory [9'd385] = 8'b10001011; 
 assign memory [9'd386] = 8'b10001000; 
 assign memory [9'd387] = 8'b10000100; 
 assign memory [9'd388] = 8'b10000000; 
 assign memory [9'd389] = 8'b01111101; 
 assign memory [9'd390] = 8'b01111001; 
 assign memory [9'd391] = 8'b01110010; 
 assign memory [9'd392] = 8'b01101011; 
 assign memory [9'd393] = 8'b01100011; 
 assign memory [9'd394] = 8'b01011100; 
 assign memory [9'd395] = 8'b01010101; 
 assign memory [9'd396] = 8'b01001110; 
 assign memory [9'd397] = 8'b01001000; 
 assign memory [9'd398] = 8'b01000001; 
 assign memory [9'd399] = 8'b00111011; 
 assign memory [9'd400] = 8'b00110101; 
 assign memory [9'd401] = 8'b00101111; 
 assign memory [9'd402] = 8'b00101001; 
 assign memory [9'd403] = 8'b00100100; 
 assign memory [9'd404] = 8'b00011111; 
 assign memory [9'd405] = 8'b00011010; 
 assign memory [9'd406] = 8'b00010110; 
 assign memory [9'd407] = 8'b00010010; 
 assign memory [9'd408] = 8'b00001110; 
 assign memory [9'd409] = 8'b00001011; 
 assign memory [9'd410] = 8'b00001000; 
 assign memory [9'd411] = 8'b00000110; 
 assign memory [9'd412] = 8'b00000100; 
 assign memory [9'd413] = 8'b00000010; 
 assign memory [9'd414] = 8'b00000001; 
 assign memory [9'd415] = 8'b00000000; 
 assign memory [9'd416] = 8'b00000000; 
 assign memory [9'd417] = 8'b00000000; 
 assign memory [9'd418] = 8'b00000000; 
 assign memory [9'd419] = 8'b00000001; 
 assign memory [9'd420] = 8'b00000010; 
 assign memory [9'd421] = 8'b00000100; 
 assign memory [9'd422] = 8'b00000110; 
 assign memory [9'd423] = 8'b00001001; 
 assign memory [9'd424] = 8'b00001100; 
 assign memory [9'd425] = 8'b00001111; 
 assign memory [9'd426] = 8'b00010001; 
 assign memory [9'd427] = 8'b00010011; 
 assign memory [9'd428] = 8'b00010101; 
 assign memory [9'd429] = 8'b00011000; 
 assign memory [9'd430] = 8'b00011010; 
 assign memory [9'd431] = 8'b00011101; 
 assign memory [9'd432] = 8'b00011111; 
 assign memory [9'd433] = 8'b00100010; 
 assign memory [9'd434] = 8'b00100101; 
 assign memory [9'd435] = 8'b00101000; 
 assign memory [9'd436] = 8'b00101011; 
 assign memory [9'd437] = 8'b00101110; 
 assign memory [9'd438] = 8'b00110010; 
 assign memory [9'd439] = 8'b00110101; 
 assign memory [9'd440] = 8'b00111000; 
 assign memory [9'd441] = 8'b00111100; 
 assign memory [9'd442] = 8'b00111111; 
 assign memory [9'd443] = 8'b01000011; 
 assign memory [9'd444] = 8'b01000111; 
 assign memory [9'd445] = 8'b01001010; 
 assign memory [9'd446] = 8'b01001110; 
 assign memory [9'd447] = 8'b01010010; 
 assign memory [9'd448] = 8'b01010110; 
 assign memory [9'd449] = 8'b01011010; 
 assign memory [9'd450] = 8'b01011110; 
 assign memory [9'd451] = 8'b01100010; 
 assign memory [9'd452] = 8'b01100110; 
 assign memory [9'd453] = 8'b01101010; 
 assign memory [9'd454] = 8'b01101110; 
 assign memory [9'd455] = 8'b01110010; 
 assign memory [9'd456] = 8'b01110110; 
 assign memory [9'd457] = 8'b01111011; 
 assign memory [9'd458] = 8'b01111111; 
 assign memory [9'd459] = 8'b10000011; 
 assign memory [9'd460] = 8'b10000111; 
 assign memory [9'd461] = 8'b10001011; 
 assign memory [9'd462] = 8'b10001111; 
 assign memory [9'd463] = 8'b10010011; 
 assign memory [9'd464] = 8'b10010111; 
 assign memory [9'd465] = 8'b10011011; 
 assign memory [9'd466] = 8'b10011111; 
 assign memory [9'd467] = 8'b10100011; 
 assign memory [9'd468] = 8'b10100111; 
 assign memory [9'd469] = 8'b10101011; 
 assign memory [9'd470] = 8'b10101111; 
 assign memory [9'd471] = 8'b10110011; 
 assign memory [9'd472] = 8'b10110111; 
 assign memory [9'd473] = 8'b10111010; 
 assign memory [9'd474] = 8'b10111110; 
 assign memory [9'd475] = 8'b11000010; 
 assign memory [9'd476] = 8'b11000101; 
 assign memory [9'd477] = 8'b11001001; 
 assign memory [9'd478] = 8'b11001100; 
 assign memory [9'd479] = 8'b11010010; 
 assign memory [9'd480] = 8'b11011001; 
 assign memory [9'd481] = 8'b11011110; 
 assign memory [9'd482] = 8'b11100100; 
 assign memory [9'd483] = 8'b11101001; 
 assign memory [9'd484] = 8'b11101101; 
 assign memory [9'd485] = 8'b11110001; 
 assign memory [9'd486] = 8'b11110101; 
 assign memory [9'd487] = 8'b11111000; 
 assign memory [9'd488] = 8'b11111010; 
 assign memory [9'd489] = 8'b11111100; 
 assign memory [9'd490] = 8'b11111110; 
 assign memory [9'd491] = 8'b11111111; 
 assign memory [9'd492] = 8'b11111111; 
 assign memory [9'd493] = 8'b11111111; 
 assign memory [9'd494] = 8'b11111111; 
 assign memory [9'd495] = 8'b11111110; 
 assign memory [9'd496] = 8'b11111100; 
 assign memory [9'd497] = 8'b11111010; 
 assign memory [9'd498] = 8'b11110111; 
 assign memory [9'd499] = 8'b11110100; 
 assign memory [9'd500] = 8'b11110000; 
 assign memory [9'd501] = 8'b11101100; 
 assign memory [9'd502] = 8'b11100111; 
 assign memory [9'd503] = 8'b11100010; 
 assign memory [9'd504] = 8'b11011101; 
 assign memory [9'd505] = 8'b11010111; 
 assign memory [9'd506] = 8'b11010001; 
 assign memory [9'd507] = 8'b11001010; 
 assign memory [9'd508] = 8'b11000011; 
 assign memory [9'd509] = 8'b10111100; 
 assign memory [9'd510] = 8'b10110100; 
 assign memory [9'd511] = 8'b10101101; 
 
endmodule


